library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY PRUEBA_VGA IS
	GENERIC(BITS:	INTEGER:=10);
	PORT(
		CLK	:	IN		STD_LOGIC;
		X		:	IN		UNSIGNED(BITS-1 DOWNTO 0);
		Y		:	IN		UNSIGNED(BITS-1 DOWNTO 0);
		RED	:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		GREEN	:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0);
		BLUE	:	OUT	STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE BEH OF PRUEBA_VGA IS
BEGIN

PROCESS (CLK)
BEGIN
	IF (RISING_EDGE(CLK)) THEN
		RED <= STD_LOGIC_VECTOR(X(4 DOWNTO 1));
		GREEN <= STD_LOGIC_VECTOR(Y(4 DOWNTO 1));
		BLUE(1 DOWNTO 0) <= STD_LOGIC_VECTOR(X(6 DOWNTO 5));
		BLUE(3 DOWNTO 2) <= STD_LOGIC_VECTOR(X(6 DOWNTO 5));
	END IF;
END PROCESS;

END ARCHITECTURE;